`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:30:57 05/11/2019 
// Design Name: 
// Module Name:    rho_tb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rho_tb(
    );
	
	reg [1599:0] state_in;
	wire [1599:0] state_out;

	assign state_in = 

	rho r(state_in, state_out)


endmodule
